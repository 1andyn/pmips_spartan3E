`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:45:55 02/21/2014 
// Design Name: 
// Module Name:    hazard_controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module hazard_controller(
    input [15:0] instruc,
	 input [2:0] opcode,
    input clock,
    output stall
    );

//Need check of Branch or Jump 
//If so, STALL

//Check for R type/ I Type




endmodule
